module L1(
    input logic end_cpu,
    output logic end_mp,

    input logic ctrl_cpu,
    output logic ctrl_mp,

    input logic status_cpu,
    output logic status_mp,

    inout logic data_cpu,
    inout logic data_mp 
);

always @(posedge clock) begin
    

end

endmodule