module L1(
    input logic end,
    output logic end,

    input logic ctrl,
    output logic ctrl,

    input logic status,
    output logic status
)