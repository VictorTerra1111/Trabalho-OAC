module mp(
    input logic end_i,
    input logic ctrl_i,

    inout logic data,
    output logic status_o
)
